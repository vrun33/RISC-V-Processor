// Wrapper conencting all the blocks

module seq_processor (
    input clk
);

    // Read from memory in initial begin


endmodule